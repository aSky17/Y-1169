//gloabl parameters for the GPU architecture

`ifndef GPU_PARAMETERS_SVH
`define GPU_PARAMETERS_SVH

package gpu_parameters;
    parameter DATA_WIDTH = 32;
    parameter OPCODE_WIDTH = 8;
    //other global p
endpackage

`endif