//gloabl parameters

`ifndef PARAMETERS_SVH
`define PARAMETERS_SVH

package parameters;
    parameter DATA_WIDTH = 32;
    parameter OPCODE_WIDTH = 8;
endpackage

`endif